`timescale 1ns / 1ps

module TWOINAND(
    );
		input A,
		input B,
		output Y
		);
		
		assign Y = A & B;

endmodule
