`timescale 1ns / 1ps

module ANDGATE(
    input A,
    input B,
    output Y
    );

	assign Y = A & B;
	
endmodule
